module overlay_creator(
    );
endmodule
